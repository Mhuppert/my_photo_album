
<h1>  <%=h @page.title %> </h1>
<br />


<%= link_to 'Edit', edit_page_path(@page) %> |
<%= link_to 'Back', pages_path %>